# Version del sistema completo 
23/02/26
V.ServerGO V0.1.1
Version = 0.1.1
