# ServerGo Version Metadata
version=0.1.2
channel=stable
release_date=2026-02-23
build=SN-F26-4
codename=Foundation
repo=https://github.com/BluePandaOpn/ServerGo
notes=Mejoras de organizacion en README/docs y menu de consola mas ordenado.
