# ServerGo Version Metadata
version=0.1.3
channel=stable
release_date=2026-02-23
build=SN-F26-5
codename=Foundation
repo=https://github.com/BluePandaOpn/ServerGo
notes=Reorganizacion completa de docs, comunidad GitHub y mejoras operativas de plataforma.
