# ServerGo Version Metadata
version=0.1.1
channel=stable
release_date=2026-02-23
build=SN-F26-2
codename=Foundation
repo=https://github.com/BluePandaOpn/ServerGo
notes=Base estable con sistema de actualizacion ZIP y docs de errores por archivo.
